library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity AxiStreamSourceMonitor_top is
generic (
    C_S_AXI_CONTROL_ADDR_WIDTH : INTEGER := 5;
    C_S_AXI_CONTROL_DATA_WIDTH : INTEGER := 32
    );
port (
    stream_clk : IN STD_LOGIC;
    s_axi_aclk : IN STD_LOGIC;
    s_axi_areset_n : IN STD_LOGIC;
    rEnable : OUT STD_LOGIC_VECTOR (0 downto 0);
    rFreerun : OUT STD_LOGIC_VECTOR (0 downto 0);
    rGeneratorSelect : OUT STD_LOGIC_VECTOR (0 downto 0);
    s_axi_control_AWVALID : IN STD_LOGIC;
    s_axi_control_AWREADY : OUT STD_LOGIC;
    s_axi_control_AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_WVALID : IN STD_LOGIC;
    s_axi_control_WREADY : OUT STD_LOGIC;
    s_axi_control_WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH/8-1 downto 0);
    s_axi_control_ARVALID : IN STD_LOGIC;
    s_axi_control_ARREADY : OUT STD_LOGIC;
    s_axi_control_ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_RVALID : OUT STD_LOGIC;
    s_axi_control_RREADY : IN STD_LOGIC;
    s_axi_control_RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    s_axi_control_BVALID : OUT STD_LOGIC;
    s_axi_control_BREADY : IN STD_LOGIC;
    s_axi_control_BRESP : OUT STD_LOGIC_VECTOR (1 downto 0)
    );
end;

architecture Behavioral of AxiStreamSourceMonitor_top is
component AxiStreamSourceMonitor is
generic (
    C_S_AXI_CONTROL_ADDR_WIDTH : INTEGER := 5;
    C_S_AXI_CONTROL_DATA_WIDTH : INTEGER := 32
);
port (
    ap_clk : IN STD_LOGIC;
    ap_rst_n : IN STD_LOGIC;
    Enable : OUT STD_LOGIC_VECTOR (0 downto 0);
    Freerun : OUT STD_LOGIC_VECTOR (0 downto 0);
    GeneratorSelect : OUT STD_LOGIC_VECTOR (0 downto 0);
    s_axi_control_AWVALID : IN STD_LOGIC;
    s_axi_control_AWREADY : OUT STD_LOGIC;
    s_axi_control_AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_WVALID : IN STD_LOGIC;
    s_axi_control_WREADY : OUT STD_LOGIC;
    s_axi_control_WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH/8-1 downto 0);
    s_axi_control_ARVALID : IN STD_LOGIC;
    s_axi_control_ARREADY : OUT STD_LOGIC;
    s_axi_control_ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_RVALID : OUT STD_LOGIC;
    s_axi_control_RREADY : IN STD_LOGIC;
    s_axi_control_RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    s_axi_control_BVALID : OUT STD_LOGIC;
    s_axi_control_BREADY : IN STD_LOGIC;
    s_axi_control_BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    interrupt : OUT STD_LOGIC
);
end component;

component HandshakeData is
generic (
    kDataWidth : natural := 8
);
port (
    InClk : in STD_LOGIC;
    OutClk : in STD_LOGIC;
    iData : in STD_LOGIC_VECTOR (kDataWidth-1 downto 0);
    oData : out STD_LOGIC_VECTOR (kDataWidth-1 downto 0);
    iPush : in STD_LOGIC;
    iRdy : out STD_LOGIC;
    oAck : in STD_LOGIC := '1';
    oValid : out STD_LOGIC;
    aiReset : in std_logic;
    aoReset : in std_logic
);
end component;

component ChangeDetectHandshake is
generic (
    kDataWidth : natural := 8
);
port (
    InClk : in STD_LOGIC;
    OutClk : in STD_LOGIC;
    iData : in STD_LOGIC_VECTOR (kDataWidth-1 downto 0);
    oData : out STD_LOGIC_VECTOR (kDataWidth-1 downto 0);
    iRdy : out STD_LOGIC;
    oValid : out STD_LOGIC;
    aiReset : in std_logic;
    aoReset : in std_logic
);
end component;

component ResetBridge is
generic (
    kPolarity : std_logic := '1'
);
port (
    aRst : in STD_LOGIC; -- asynchronous reset; active-high, if kPolarity=1
    OutClk : in STD_LOGIC;
    oRst : out STD_LOGIC
);
end component;

-- HLS interrupt flag
signal lInterrupt : STD_LOGIC;

-- Reset signals for each clock domain
signal rRst_n : STD_LOGIC;
signal rRst : STD_LOGIC;
signal lRst_n : STD_LOGIC;
signal lRst : STD_LOGIC;

-- Internal signals for ports
signal lEnable : STD_LOGIC_VECTOR (0 downto 0);
signal rEnableInt : STD_LOGIC_VECTOR (0 downto 0);
signal lFreerun : STD_LOGIC_VECTOR (0 downto 0);
signal rFreerunInt : STD_LOGIC_VECTOR (0 downto 0);
signal lGeneratorSelect : STD_LOGIC_VECTOR (0 downto 0);
signal rGeneratorSelectInt : STD_LOGIC_VECTOR (0 downto 0);


begin

--- Instantiate HLS register file core

AxiStreamSourceMonitor_inst: AxiStreamSourceMonitor port map(
    ap_clk => s_axi_aclk,
    ap_rst_n => s_axi_areset_n,
    Enable => lEnable,
    Freerun => lFreerun,
    GeneratorSelect => lGeneratorSelect,
    s_axi_control_AWVALID => s_axi_control_AWVALID,
    s_axi_control_AWREADY => s_axi_control_AWREADY,
    s_axi_control_AWADDR => s_axi_control_AWADDR,
    s_axi_control_WVALID => s_axi_control_WVALID,
    s_axi_control_WREADY => s_axi_control_WREADY,
    s_axi_control_WDATA => s_axi_control_WDATA,
    s_axi_control_WSTRB => s_axi_control_WSTRB,
    s_axi_control_ARVALID => s_axi_control_ARVALID,
    s_axi_control_ARREADY => s_axi_control_ARREADY,
    s_axi_control_ARADDR => s_axi_control_ARADDR,
    s_axi_control_RVALID => s_axi_control_RVALID,
    s_axi_control_RREADY => s_axi_control_RREADY,
    s_axi_control_RDATA => s_axi_control_RDATA,
    s_axi_control_RRESP => s_axi_control_RRESP,
    s_axi_control_BVALID => s_axi_control_BVALID,
    s_axi_control_BREADY => s_axi_control_BREADY,
    s_axi_control_BRESP => s_axi_control_BRESP,
    interrupt => lInterrupt
);

--- Create synchronous resets for each clock

s_axi_aclk_to_stream_clk_rst: ResetBridge generic map(
    kPolarity => '0'
)
port map (
    aRst => s_axi_areset_n,
    outClk => stream_clk,
    oRst => rRst_n
);
rRst <= not rRst_n;
lRst_n <= s_axi_areset_n;
lRst <= not s_axi_areset_n;

--- Map external output ports to internal signals
rEnable <= rEnableInt;
rFreerun <= rFreerunInt;
rGeneratorSelect <= rGeneratorSelectInt;

--- Instantiate handshake clock domain crossing modules
-- Handshake CDC for Enable from s_axi_aclk to stream_clk
--- trigger handshake on HLS interrupt
Enable_from_s_axi_aclk_to_stream_clk_InstHandshake: HandshakeData 
generic map (
    kDataWidth => 1
)
port map(
    InClk => s_axi_aclk,
    OutClk => stream_clk,
    iData => lEnable,
    oData => rEnableInt,
    iPush => lInterrupt,
    iRdy => open,
    oAck => '1',
    oValid => open,
    aiReset => lRst,
    aoReset => rRst
);
-- Handshake CDC for Freerun from s_axi_aclk to stream_clk
--- trigger handshake on HLS interrupt
Freerun_from_s_axi_aclk_to_stream_clk_InstHandshake: HandshakeData 
generic map (
    kDataWidth => 1
)
port map(
    InClk => s_axi_aclk,
    OutClk => stream_clk,
    iData => lFreerun,
    oData => rFreerunInt,
    iPush => lInterrupt,
    iRdy => open,
    oAck => '1',
    oValid => open,
    aiReset => lRst,
    aoReset => rRst
);
-- Handshake CDC for GeneratorSelect from s_axi_aclk to stream_clk
--- trigger handshake on HLS interrupt
GeneratorSelect_from_s_axi_aclk_to_stream_clk_InstHandshake: HandshakeData 
generic map (
    kDataWidth => 1
)
port map(
    InClk => s_axi_aclk,
    OutClk => stream_clk,
    iData => lGeneratorSelect,
    oData => rGeneratorSelectInt,
    iPush => lInterrupt,
    iRdy => open,
    oAck => '1',
    oValid => open,
    aiReset => lRst,
    aoReset => rRst
);

end Behavioral;
